LIBRARY IEEE;
USE IEEE.std_logic_1164.all;

ENTITY mux8x1 IS 
	Generic ( n : Integer:=16);
	PORT ( in0,in1,in2,in3,in4,in5,in6,in7 : IN std_logic_vector (n-1 DOWNTO 0);
			sel : IN  std_logic_vector (1 DOWNTO 0);
			out1 : OUT std_logic_vector (n-1 DOWNTO 0));
END entity;


ARCHITECTURE when_else_mux2 OF mux8x1 is
	BEGIN
		
  out1 <= 	in0 when sel = "000"
	else	in1 when sel = "001"
	else	in2 when sel = "010"
	else 	in3  when sel = "011"
	else in4 when sel = "100"
	else in5 when sel = "101"
	else in6 when sel = "110"
	else in7;
	
END when_else_mux2;

