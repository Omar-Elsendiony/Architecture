Library ieee;
Use ieee.std_logic_1164.all;
Package mine is

Constant zeroFlag : integer :=0;
Constant carryFlag : integer :=1;
Constant negativeFlag : integer :=2;

--Constant RegWrite : integer :=12;
--Constant MemWrite : integer :=12;
--Constant MemRead : integer :=12;
--Constant ALUFn : integer :=12;
--Constant RegInSrc : integer :=12;
--Constant SPEn : integer :=12;
--Constant SPStatus : integer :=12;

End mine;